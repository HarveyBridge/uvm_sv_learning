
module test_top;
	$display("hello 123");
endmodule
