
module test_top;
	$display("hello");
endmodule
